module plugin

@[if debug]
fn debug(s string) {
	eprintln(s)
}

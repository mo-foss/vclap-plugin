module vclap

@[if debug]
fn debug(s string) {
	eprintln(s)
}
